library ieee;
use ieee.std_logic_1164.all;
entity hex_to_sseg is
	port(
		clk    : in  std_logic;
		reset  : in  std_logic;
		hex    : in  std_logic_vector(3 downto 0);
		dp     : in  std_logic;
		sseg_o : out std_logic_vector(7 downto 0)
	);
end hex_to_sseg;

architecture arch of hex_to_sseg is
	signal sseg : std_logic_vector(7 downto 0);
begin

	process(clk, reset, sseg)
	begin
		if (reset = '1') then
			sseg_o <= (others => '1');
		elsif rising_edge(clk) then
			sseg_o <= not sseg;
		end if;
	end process;

	with hex select sseg(6 downto 0) <=
		"0000001" when "0000",
		"1001111" when "0001",
		"0010010" when "0010",
		"0000110" when "0011",
		"1001100" when "0100",
		"0100100" when "0101",
		"0100000" when "0110",
		"0001111" when "0111",
		"0000000" when "1000",
		"0000100" when "1001",
		"0001000" when "1010",         --a
		"1100000" when "1011",         --b
		"0110001" when "1100",         --c
		"1000010" when "1101",         --d
		"0110000" when "1110",         --e
		"0111000" when others;         --f
		
	-- decimal point
	sseg(7) <= dp;
end arch;
