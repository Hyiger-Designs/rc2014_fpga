cpu_data_inst : cpu_data PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataio	 => dataio_sig,
		dataout	 => dataout_sig
	);
