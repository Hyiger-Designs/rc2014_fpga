data_bus_inst : data_bus PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataio	 => dataio_sig,
		dataout	 => dataout_sig
	);
