library IEEE;
use IEEE.STD_LOGIC_1164.all;

package user_types is

	type sseg is array (0 to 5) of std_logic_vector(7 downto 0);

end user_types;

package body user_types is

end user_types;
